module TwiddleX ( 
	input logic [15:0] Xr,
    input logic [15:0] Yr,
	input logic  [15:0] Xi,
    input logic  [15:0] Yi,
    input logic clk,
    output logic overflow,       
    output logic  [31:0] Outr,
    output logic  [31:0] Outi
);

endmodule